module font_rom_state(input [5:0] addr, 
					output [15:0] data);
					
					
parameter ADDR_WIDTH = 6;
parameter DATA_WIDTH = 16;
logic [ADDR_WIDTH-1:0] addr_reg;
assign data = ROM[addr];

parameter [0:2**ADDR_WIDTH-1][DATA_WIDTH-1:0] ROM = {
	//x0C
	16'b0000000000000000,//1
	16'b0110000000000110,//0//over, cross, X
	16'b0111000000001110,//2
	16'b0011100000011100,//3
	16'b0001110000111000,//4
	16'b0000111001110000,//5
	16'b0000011111100000,//6
	16'b0000001111000000,//7
	16'b0000000110000000,//16
	16'b0000001111000000,//9
	16'b0000011111100000,//1
	16'b0000111001110000,//1
	16'b0001110000111000,//1
	16'b0011100000011100,//1
	16'b0111000000001110,//1
	16'b0110000000000110,//1
	//x0A
	//x0B
	16'b0000000000000000,//1
	16'b0111110000111110,//1
	16'b0111110000111110,//1
	16'b0111110000111110,//1
	16'b0111110000111110,//1
	16'b0111110000111110,//1
	16'b0111110000111110,//1
	16'b0111110000111110,//1
	16'b0111110000111110,//1
	16'b0111110000111110,//1
	16'b0111110000111110,//1
	16'b0111110000111110,//1
	16'b0111110000111110,//1
	16'b0111110000111110,//1
	16'b0111110000111110,//1
	16'b0000000000000000,//1
	
	
	16'b0000000000000000,//1
	16'b0100000000000000,//1
	16'b0111000000000000,//1
	16'b0111110000000000,//1
	16'b0111111110000000,//1
	16'b0111111111000000,//1
	16'b0111111111110000,//1
	16'b0111111111111100,//1
	16'b0111111111111110,//1
	16'b0111111111111100,//1
	16'b0111111111110000,//1
	16'b0111111111000000,//1
	16'b0111111100000000,//1
	16'b0111110000000000,//1
	16'b0111000000000000,//1
	16'b0100000000000000,//1
	
	
		//x0C
	16'b0000000000000000,//1
	16'b1110000000000111,//0//over, cross, X
	16'b0111000000001110,//2
	16'b0011100000011100,//3
	16'b0001110000111000,//4
	16'b0000111001110000,//5
	16'b0000011111100000,//6
	16'b0000001111000000,//7
	16'b000000011000000,//16
	16'b0000001111000000,//9
	16'b0000011111100000,//1
	16'b0000111001110000,//1
	16'b0001110000111000,//1
	16'b0011100000011100,//1
	16'b0111000000001110,//1
	16'b1110000000000111//1
	
	
	
	
	
	
};

endmodule
