module font_rom_num(input [6:0] addr, 
					output [7:0] data);
					
					
parameter ADDR_WIDTH = 7;
parameter DATA_WIDTH = 8;
logic [ADDR_WIDTH-1:0] addr_reg;
assign data = ROM[addr];

parameter [0:2**ADDR_WIDTH-1][DATA_WIDTH-1:0] ROM = {
	8'b00000000,//0//zero
	8'b00111100,//1
	8'b01111110,//2
	8'b01100110,//3
	8'b01100110,//4
	8'b01100110,//5
	8'b01100110,//6
	8'b01111110,//7
	8'b00111100,//8
	8'b00000000,//9
	//x03
	8'b00000000,//0//one
	8'b00011000,//1
	8'b00111000,//2
	8'b01111000,//3
	8'b00011000,//4
	8'b00011000,//5
	8'b00011000,//6
	8'b00011000,//7
	8'b01111110,//8
	8'b00000000,//9
	//x01
	8'b00000000,//0//two
	8'b01111110,//1
	8'b01111110,//2
	8'b00000110,//3
	8'b01111110,//4
	8'b01111110,//5
	8'b01100000,//6
	8'b01111110,//7
	8'b01111110,//8
	8'b00000000,//9
	//x01
	8'b00000000,//0//three
	8'b01111110,//1
	8'b01111110,//2
	8'b00000110,//3
	8'b01111110,//4
	8'b01111110,//5
	8'b00000110,//6
	8'b01111110,//7
	8'b01111110,//8
	8'b00000000,//9
	//x01
	8'b00000000,//0//four
	8'b01100110,//1
	8'b01100110,//2
	8'b01100110,//3
	8'b01111110,//4
	8'b00000110,//5
	8'b00000110,//6
	8'b00000110,//7
	8'b00000110,//8
	8'b00000000,//9
	//x01
	8'b00000000,//0//five
	8'b01111110,//1
	8'b01111110,//2
	8'b01100000,//3
	8'b01111110,//4
	8'b01111110,//5
	8'b00000110,//6
	8'b01111110,//7
	8'b01111110,//8
	8'b00000000,//9
	//x01
	8'b00000000,//0//six
	8'b01111110,//1
	8'b01111110,//2
	8'b01100000,//3
	8'b01111110,//4
	8'b01111110,//5
	8'b01100110,//6
	8'b01111110,//7
	8'b01111110,//8
	8'b00000000,//9
	//x01
	8'b00000000,//0//seven
	8'b01111110,//1
	8'b01111110,//2
	8'b00000110,//3
	8'b00000110,//4
	8'b00000110,//5
	8'b00000110,//6
	8'b00000110,//7
	8'b00000110,//8
	8'b00000000,//9
	//x01
	8'b00000000,//0//eight
	8'b01111110,//1
	8'b01111110,//2
	8'b01100110,//3
	8'b01111110,//4
	8'b01111110,//5
	8'b01100110,//6
	8'b01111110,//7
	8'b01111110,//8
	8'b00000000,//9
	//x01
	8'b00000000,//0//nine
	8'b01111110,//1
	8'b01111110,//2
	8'b01100110,//3
	8'b01111110,//4
	8'b01111110,//5
	8'b00000110,//6
	8'b01111110,//7
	8'b01111110,//8
	8'b00000000,//9
	
	//trash
	8'b00000000,//0//zero
	8'b00111100,//1
	8'b01111110,//2
	8'b01100110,//3
	8'b01100110,//4
	8'b01100110,//5
	8'b01100110,//6
	8'b01111110,//7
	8'b00111100,//8
	8'b00000000,//9
	//x03
	8'b00000000,//0//one
	8'b00011000,//1
	8'b00111000,//2
	8'b01111000,//3
	8'b00011000,//4
	8'b00011000,//5
	8'b00011000,//6
	8'b00011000,//7
	8'b01111110,//8
	8'b00000000,//9
	//x01
	8'b00000000,//0//two
	8'b01111110,//1
	8'b01111110,//2
	8'b00000110,//3
	8'b01111110,//4
	8'b01111110,//5
	8'b01100000,//6
	8'b01111110//7
};

endmodule
