module font_rom_enter(input [7:0] addr, 
					output [7:0] data);
					
					
parameter ADDR_WIDTH =8;
parameter DATA_WIDTH = 8;
logic [ADDR_WIDTH-1:0] addr_reg;
assign data = ROM[addr];

parameter [0:2**ADDR_WIDTH-1][DATA_WIDTH-1:0] ROM = {
	//x01
	8'b00000000,//0//P
	8'b01111110,//2
	8'b01111110,//31
	8'b01100110,//4
	8'b01111110,//5
	8'b01111110,//6
	8'b01100000,//7
	8'b01100000,//8
	8'b01100000,//9
	8'b00000000,//1
	//x01
	8'b00000000,//0//R
	8'b01111110,//1
	8'b01111110,//2
	8'b01100110,//3
	8'b01111110,//4
	8'b01111000,//5
	8'b01101100,//6
	8'b01100110,//7
	8'b01100010,//8
	8'b00000000,//9
	//x02
	8'b00000000,//0//E
	8'b01111110,//1
	8'b01111110,//2
	8'b01100000,//3
	8'b01111110,//4
	8'b01111110,//5
	8'b01100000,//6
	8'b01111110,//7
	8'b01111110,//8
	8'b00000000,//9
	//x03
	8'b00000000,//0//S
	8'b01111110,//1
	8'b01111110,//2
	8'b01100000,//3
	8'b01111110,//4
	8'b01111110,//5
	8'b00000110,//6
	8'b01111110,//7
	8'b01111110,//8
	8'b00000000,//9
	//x04
	8'b00000000,//0//S
	8'b01111110,//1
	8'b01111110,//2
	8'b01100000,//3
	8'b01111110,//4
	8'b01111110,//5
	8'b00000110,//6
	8'b01111110,//7
	8'b01111110,//8
	8'b00000000,//9
	//x06
	//x00
	8'b00000000,//0//space
	8'b00000000,//1
	8'b00000000,//2
	8'b00000000,//3
	8'b00000000,//4
	8'b00000000,//5
	8'b00000000,//6
	8'b00000000,//7
	8'b00000000,//8
	8'b00000000,//9
	//x01
	8'b00000000,//0//E
	8'b01111110,//1
	8'b01111110,//2
	8'b01100000,//3
	8'b01111110,//4
	8'b01111110,//5
	8'b01100000,//6
	8'b01111110,//7
	8'b01111110,//8
	8'b00000000,//9
	//x03
	8'b00000000,//0//N
	8'b01111110,//2
	8'b01111110,//3
	8'b01100110,//4
	8'b01100110,//5
	8'b01100110,//6
	8'b01100110,//7
	8'b01100110,//8
	8'b01100110,//9
	8'b00000000,//1
	//x08
	8'b00000000,//0//T
	8'b01111110,//1
	8'b01111110,//2
	8'b00011000,//3
	8'b00011000,//4
	8'b00011000,//5
	8'b00011000,//6
	8'b00011000,//7
	8'b00011000,//8
	8'b00000000,//9
	//x02
	8'b00000000,//0//E
	8'b01111110,//1
	8'b01111110,//2
	8'b01100000,//3
	8'b01111110,//4
	8'b01111110,//5
	8'b01100000,//6
	8'b01111110,//7
	8'b01111110,//8
	8'b00000000,//9
	//x03
	8'b00000000,//0//R
	8'b01111110,//1
	8'b01111110,//2
	8'b01100110,//3
	8'b01111110,//4
	8'b01111000,//5
	8'b01101100,//6
	8'b01100110,//7
	8'b01100010,//8
	8'b00000000,//9
	//x04
	8'b00000000,//0//space
	8'b00000000,//1
	8'b00000000,//2
	8'b00000000,//3
	8'b00000000,//4
	8'b00000000,//5
	8'b00000000,//6
	8'b00000000,//7
	8'b00000000,//8
	8'b00000000,//9
	//x01
	8'b00000000,//0//T
	8'b01111110,//1
	8'b01111110,//2
	8'b00011000,//3
	8'b00011000,//4
	8'b00011000,//5
	8'b00011000,//6
	8'b00011000,//7
	8'b00011000,//8
	8'b00000000,//9
	//x02
	8'b00000000,//0//O
	8'b01111110,//1
	8'b01111110,//2
	8'b01100110,//3
	8'b01100110,//4
	8'b01100110,//5
	8'b01100110,//6
	8'b01111110,//7
	8'b01111110,//8
	8'b00000000,//9
	
	8'b00000000,//0//space
	8'b00000000,//1
	8'b00000000,//2
	8'b00000000,//3
	8'b00000000,//4
	8'b00000000,//5
	8'b00000000,//6
	8'b00000000,//7
	8'b00000000,//8
	8'b00000000,//9
	//x01
	8'b00000000,//0//B
	8'b01111100,//1
	8'b01111110,//2
	8'b01100110,//3
	8'b01111110,//4
	8'b01111110,//5
	8'b01100110,//6
	8'b01111110,//7
	8'b01111100,//8
	8'b00000000,//9
	
	8'b00000000,//0//E
	8'b01111110,//1
	8'b01111110,//2
	8'b01100000,//3
	8'b01111110,//4
	8'b01111110,//5
	8'b01100000,//6
	8'b01111110,//7
	8'b01111110,//8
	8'b00000000,//9
	
	8'b00000000,//0//G
	8'b01111110,//1
	8'b01111110,//2
	8'b01100000,//3
	8'b01101110,//4
	8'b01101110,//5
	8'b01100110,//6
	8'b01111110,//7
	8'b01111110,//8
	8'b00000000,//9
	
	//x09
	8'b00000000,//0//I
	8'b01111110,//1
	8'b01111110,//2
	8'b00011000,//3
	8'b00011000,//4
	8'b00011000,//5
	8'b00011000,//6
	8'b01111110,//7
	8'b01111110,//8
	8'b00000000,//9
	//x05
	8'b00000000,//0//N
	8'b01111110,//2
	8'b01111110,//3
	8'b01100110,//4
	8'b01100110,//5
	8'b01100110,//6
	8'b01100110,//7
	8'b01100110,//8
	8'b01100110,//9
	8'b00000000,//1
	//x08	
	//trash
	8'b00000000,//0//N
	8'b01111110,//2
	8'b01111110,//3
	8'b01100110,//4
	8'b01100110,//5
	8'b01100110,//6
	8'b01100110,//7
	8'b01100110,//8
	8'b01100110,//9
	8'b00000000,//1
	8'b00000000,//0//N
	8'b01111110,//2
	8'b01111110,//3
	8'b01100110,//4
	8'b01100110,//5
	8'b01100110,//6
	8'b01100110,//7
	8'b01100110,//8
	8'b01100110,//9
	8'b00000000,//1
	8'b00000000,//0//N
	8'b01111110,//2
	8'b01111110,//3
	8'b01100110,//4
	8'b01100110,//5
	8'b01100110,//6
	8'b01100110,//7
	8'b01100110,//8
	8'b01100110,//9
	8'b00000000,//1
	8'b00000000,//0//N
	8'b01111110,//2
	8'b01111110,//3
	8'b01100110,//4
	8'b01100110,//5
	8'b01100110,//6
	8'b01100110,//7
	8'b01100110,//8
	8'b01100110,//9
	8'b00000000,//1
	8'b00000000,//0//N
	8'b01111110,//2
	8'b01111110,//3
	8'b01100110,//4
	8'b01100110,//5
	8'b01100110,//6
	8'b01100110,//7
	8'b01100110,//8
	8'b01100110,//9
	8'b00000000,//1
	8'b00000000,//0//N
	8'b01111110,//2
	8'b01111110,//3
	8'b01100110,//4
	8'b01100110,//5
	8'b01100110//6
};

endmodule
